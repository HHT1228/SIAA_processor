module InstrROM #(parameter D=8)(
  input       [D-1:0] addr,    // prog_ctr	  address pointer
  output logic [8:0] readData);

  logic[8:0] memory[2**D];
  initial begin							    // load the program
		$readmemb("F:/UCSD/WI23/CSE 141L/SIAA/Program1/mach_code.txt", memory);
	end

  always_comb  readData = memory[addr];

endmodule

